package pkg;


//import uvm_pkg.sv
	import uvm_pkg::*;
//include uvm_macros.sv
	`include "uvm_macros.svh"
//`include "tb_defs.sv"
`include "src_xtn.sv"
`include "src_agt_cfg.sv"
`include "dst_agt_cfg.sv"
`include "env_config.sv"
`include "src_drv.sv"
`include "src_mon.sv"
`include "src_sequencer.sv"
`include "src_agent.sv"
`include "src_agt_top.sv"
`include "src_seq.sv"

`include "dst_xtn.sv"
`include "dst_mon.sv"
`include "dst_sequencer.sv"
`include "dst_sequence.sv"
`include "dst_drv.sv"
`include "dst_agent.sv"
`include "dst_agent_top.sv"

`include "router_virtual_sequencer.sv"
`include "virtual_seq.sv"
`include "scoreboard.sv"

`include "router_env.sv"


`include "test.sv"
endpackage
